`timescale 1ns / 1ns
module test;

    reg [7:0] num;      
    wire result;         

    is_even testing_module (
        .num(num),
        .result(result)
    );

    initial begin
        num = 8'd0;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd1;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd2;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd3;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd4;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd5;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd6;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd7;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd8;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd9;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd10;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd11;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd12;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd13;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd14;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd15;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd16;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd17;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd18;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd19;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd20;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd21;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd22;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd23;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd24;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd25;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd26;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd27;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd28;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd29;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd30;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd31;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd32;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd33;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd34;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd35;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd36;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd37;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd38;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd39;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd40;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd41;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd42;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd43;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd44;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd45;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd46;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd47;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd48;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd49;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd50;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd51;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd52;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd53;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd54;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd55;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd56;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd57;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd58;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd59;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd60;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd61;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd62;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd63;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd64;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd65;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd66;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd67;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd68;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd69;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd70;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd71;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd72;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd73;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd74;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd75;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd76;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd77;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd78;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd79;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd80;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd81;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd82;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd83;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd84;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd85;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd86;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd87;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd88;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd89;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd90;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd91;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd92;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd93;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd94;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd95;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd96;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd97;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd98;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd99;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd100;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd101;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd102;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd103;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd104;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd105;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd106;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd107;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd108;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd109;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd110;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd111;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd112;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd113;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd114;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd115;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd116;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd117;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd118;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd119;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd120;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd121;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd122;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd123;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd124;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd125;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd126;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd127;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd128;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd129;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd130;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd131;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd132;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd133;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd134;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd135;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd136;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd137;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd138;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd139;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd140;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd141;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd142;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd143;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd144;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd145;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd146;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd147;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd148;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd149;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd150;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd151;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd152;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd153;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd154;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd155;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd156;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd157;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd158;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd159;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd160;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd161;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd162;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd163;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd164;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd165;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd166;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd167;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd168;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd169;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd170;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd171;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd172;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd173;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd174;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd175;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd176;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd177;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd178;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd179;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd180;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd181;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd182;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd183;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd184;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd185;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd186;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd187;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd188;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd189;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd190;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd191;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd192;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd193;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd194;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd195;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd196;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd197;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd198;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd199;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd200;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd201;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd202;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd203;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd204;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd205;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd206;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd207;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd208;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd209;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd210;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd211;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd212;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd213;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd214;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd215;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd216;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd217;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd218;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd219;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd220;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd221;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd222;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd223;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd224;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd225;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd226;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd227;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd228;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd229;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd230;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd231;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd232;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd233;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd234;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd235;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd236;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd237;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd238;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd239;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd240;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd241;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd242;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd243;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd244;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd245;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd246;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd247;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd248;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd249;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd250;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd251;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd252;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd253;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd254;  #1000000000; $display("%d \t %b", num, result);
        num = 8'd255;  #1000000000; $display("%d \t %b", num, result);

        $stop;
    end
endmodule
